`timescale 1ns / 1ps 

module EFCDT (Va,Vb,Vc,Ia,Ib,Ic,cls);

parameter N = 'd8;
parameter C = 'd3;
input logic[N-1:0] Va,Vb,Vc,Ia,Ib,Ic;
output logic [C-1:0] cls;

logic ns0,ns1,ns2,ns3,ns4,ns7,ns10,ns11,ns14,ns17,ns18,ns19,ns23,ns24,ns27,ns30,ns31,ns32,ns33,ns36,ns39,ns40,ns43,ns46,ns47,ns50;
parameter logic[N-1:0] t0 = 8'd137;
parameter logic[N-1:0] t1 = 8'd136;
parameter logic[N-1:0] t2 = 8'd117;
parameter logic[N-1:0] t3 = 8'd134;
parameter logic[N-1:0] t4 = 8'd114;
parameter logic[N-1:0] t7 = 8'd122;
parameter logic[N-1:0] t10 = 8'd143;
parameter logic[N-1:0] t11 = 8'd123;
parameter logic[N-1:0] t14 = 8'd112;
parameter logic[N-1:0] t17 = 8'd120;
parameter logic[N-1:0] t18 = 8'd231;
parameter logic[N-1:0] t19 = 8'd159;
parameter logic[N-1:0] t23 = 8'd122;
parameter logic[N-1:0] t24 = 8'd172;
parameter logic[N-1:0] t27 = 8'd140;
parameter logic[N-1:0] t30 = 8'd138;
parameter logic[N-1:0] t31 = 8'd120;
parameter logic[N-1:0] t32 = 8'd120;
parameter logic[N-1:0] t33 = 8'd134;
parameter logic[N-1:0] t36 = 8'd161;
parameter logic[N-1:0] t39 = 8'd128;
parameter logic[N-1:0] t40 = 8'd122;
parameter logic[N-1:0] t43 = 8'd89;
parameter logic[N-1:0] t46 = 8'd133;
parameter logic[N-1:0] t47 = 8'd125;
parameter logic[N-1:0] t50 = 8'd184;

assign ns0 = (Ic < t0)? 1:0;
assign ns1 = (Ia < t1)? 1:0;
assign ns2 = (Ia < t2)? 1:0;
assign ns3 = (Ib < t3)? 1:0;
assign ns4 = (Ib < t4)? 1:0;
assign ns7 = (Ic < t7)? 1:0;
assign ns10 = (Ib < t10)? 1:0;
assign ns11 = (Ib < t11)? 1:0;
assign ns14 = (Vb < t14)? 1:0;
assign ns17 = (Ic < t17)? 1:0;
assign ns18 = (Ib < t18)? 1:0;
assign ns19 = (Vc < t19)? 1:0;
assign ns23 = (Ib < t23)? 1:0;
assign ns24 = (Vc < t24)? 1:0;
assign ns27 = (Ib < t27)? 1:0;
assign ns30 = (Vc < t30)? 1:0;
assign ns31 = (Vc < t31)? 1:0;
assign ns32 = (Ib < t32)? 1:0;
assign ns33 = (Vb < t33)? 1:0;
assign ns36 = (Ib < t36)? 1:0;
assign ns39 = (Va < t39)? 1:0;
assign ns40 = (Va < t40)? 1:0;
assign ns43 = (Ia < t43)? 1:0;
assign ns46 = (Vb < t46)? 1:0;
assign ns47 = (Ib < t47)? 1:0;
assign ns50 = (Ib < t50)? 1:0;

always_comb
begin
    casex({ns0,ns1,ns2,ns3,ns4,ns7,ns10,ns11,ns14,ns17,ns18,ns19,ns23,ns24,ns27,ns30,ns31,ns32,ns33,ns36,ns39,ns40,ns43,ns46,ns47,ns50})
		26'b11111?????????????????????: cls = 'd2;
		26'b11110?????????????????????: cls = 'd1;
		26'b1110?1????????????????????: cls = 'd5;
		26'b1110?0????????????????????: cls = 'd2;
		26'b110???11??????????????????: cls = 'd2;
		26'b110???10??????????????????: cls = 'd0;
		26'b110???0?1?????????????????: cls = 'd2;
		26'b110???0?0?????????????????: cls = 'd4;
		26'b10???????111??????????????: cls = 'd3;
		26'b10???????110??????????????: cls = 'd5;
		26'b10???????10???????????????: cls = 'd3;
		26'b10???????0??11????????????: cls = 'd2;
		26'b10???????0??10????????????: cls = 'd5;
		26'b10???????0??0?1???????????: cls = 'd1;
		26'b10???????0??0?0???????????: cls = 'd2;
		26'b0??????????????1111???????: cls = 'd4;
		26'b0??????????????1110???????: cls = 'd4;
		26'b0??????????????110?1??????: cls = 'd3;
		26'b0??????????????110?0??????: cls = 'd3;
		26'b0??????????????10???11????: cls = 'd3;
		26'b0??????????????10???10????: cls = 'd3;
		26'b0??????????????10???0?1???: cls = 'd5;
		26'b0??????????????10???0?0???: cls = 'd4;
		26'b0??????????????0???????11?: cls = 'd4;
		26'b0??????????????0???????10?: cls = 'd4;
		26'b0??????????????0???????0?1: cls = 'd3;
		26'b0??????????????0???????0?0: cls = 'd5;
		default: cls = '0;
	endcase
end

endmodule
